-- package to print traces of cmd executions
-- TODO