library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.conversions_pack.all;
use work.cpu_defs_pack.all;

package instr_encode_pack is

end instr_encode_pack;

package body instr_encode_pack is

end instr_encode_pack;